library verilog;
use verilog.vl_types.all;
entity id_sv_unit is
end id_sv_unit;
