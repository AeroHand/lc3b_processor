library verilog;
use verilog.vl_types.all;
entity adjz_sv_unit is
end adjz_sv_unit;
