library verilog;
use verilog.vl_types.all;
entity wb_sv_unit is
end wb_sv_unit;
