library verilog;
use verilog.vl_types.all;
entity ifetch_sv_unit is
end ifetch_sv_unit;
