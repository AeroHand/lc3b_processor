library verilog;
use verilog.vl_types.all;
entity cache2_sv_unit is
end cache2_sv_unit;
