library verilog;
use verilog.vl_types.all;
entity forward_unit_sv_unit is
end forward_unit_sv_unit;
