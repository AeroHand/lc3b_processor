library verilog;
use verilog.vl_types.all;
entity write_calc_sv_unit is
end write_calc_sv_unit;
