library verilog;
use verilog.vl_types.all;
entity tagcomp_sv_unit is
end tagcomp_sv_unit;
