library verilog;
use verilog.vl_types.all;
entity off_addr_calc_sv_unit is
end off_addr_calc_sv_unit;
