library verilog;
use verilog.vl_types.all;
entity cache_datapath_2_sv_unit is
end cache_datapath_2_sv_unit;
