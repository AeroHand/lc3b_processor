library verilog;
use verilog.vl_types.all;
entity ex_sv_unit is
end ex_sv_unit;
