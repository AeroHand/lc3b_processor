library verilog;
use verilog.vl_types.all;
entity nzp_comparator_sv_unit is
end nzp_comparator_sv_unit;
